module yima(Q,Q1,Q2);
input [7:0]Q;
output reg [6:0]Q1;
output reg [6:0]Q2;
reg [3:0]q1;
reg [3:0]q2;
always @ (Q)
begin 
q1[0]=Q[0];
q1[1]=Q[1];
q1[2]=Q[2];
q1[3]=Q[3];
q2[0]=Q[4];
q2[1]=Q[5];
q2[2]=Q[6];
q2[3]=Q[7];
Q1=7'b0000000;
Q2=7'b0000000;
case(q1)
4'b0000:Q1=7'b0111111;
4'b0001:Q1=7'b0000110;
4'b0010:Q1=7'b1011011;
4'b0011:Q1=7'b1001111;
4'b0100:Q1=7'b1100110;
4'b0101:Q1=7'b1101101;
4'b0110:Q1=7'b1111100;
4'b0111:Q1=7'b0000111;
4'b1000:Q1=7'b1111111;
4'b1001:Q1=7'b1100111;
default:Q1=7'b0000000;
endcase
case(q2)
4'b0000:Q2=7'b0111111;
4'b0001:Q2=7'b0000110;
4'b0010:Q2=7'b1011011;
4'b0011:Q2=7'b1001111;
4'b0100:Q2=7'b1100110;
4'b0101:Q2=7'b1101101;
4'b0110:Q2=7'b1111100;
4'b0111:Q2=7'b0000111;
4'b1000:Q2=7'b1111111;
4'b1001:Q2=7'b1100111;
default:Q2=7'b0000000;
endcase
end 
endmodule 


